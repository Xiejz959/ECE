LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MUX4bit4to1 IS
	PORT 
	(
        U   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);  
        V   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);  
        W   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);  
        X   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);  
        S   : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);  -- S1=S[1], S0=S[0]
        M   : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)   
    );

END MUX4bit4to1;

ARCHITECTURE comb OF MUX4bit4to1 IS
BEGIN
	WITH S SELECT
	M <= U WHEN "00", --00
		  V WHEN "10", --10
		  W WHEN "01", --01
		  X WHEN OTHERS;

END comb;
